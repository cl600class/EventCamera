// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// PROGRAM		"Quartus II 64-Bit"
// VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
// CREATED		"Thu May 30 01:31:16 2019"



module asymc(
	I0,
	I1,
	Q
);


input wire	I0;
input wire	I1;
output wire	Q;

wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;

assign	Q = SYNTHESIZED_WIRE_0;




or_2	b2v_inst(
	.i1(SYNTHESIZED_WIRE_0),
	.i2(I1),
	.o1(SYNTHESIZED_WIRE_1));


and_2	b2v_inst5(
	.i1(SYNTHESIZED_WIRE_1),
	.i2(I0),
	.o1(SYNTHESIZED_WIRE_0));


endmodule
